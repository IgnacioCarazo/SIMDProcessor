module decoder #(parameter N=24, parameter registerSize = 32)
                 (input logic [N-1:0] instruction,  // Instrucción de N bits
                  output logic MemoryWrite,          // Control para escribir en memoria
                  output logic [1:0] WriteRegFrom,   // Indica de dónde provienen los datos que vamos a escribir en el registro
                  output logic [3:0] RegToWrite,     // Registro donde se escriben los datos
                  output logic [registerSize - 1:0] Immediate, // Valor inmediato extraído de la instrucción
                  output logic writeMemFrom,         // Control que indica si los datos a escribir en memoria provienen de la instrucción.
                  output logic RegWriteEnSc,         // Habilitación de escritura en registro escalar
                  output logic RegWriteEnVec,        // Habilitación de escritura en registro vectorial
                  output logic [2:0] PcWriteEn,      // Control para escribir en el PC
                  output logic OverWriteNz,          // Bandera para sobrescribir NZ (flags de condición)
                  output logic [2:0] AluOpCode       // Código de operación para la ALU
);

    logic memoryInstruction, regWriteEn, preliminar_write_reg_from_1;
    logic jump_instruction;
		
    assign jump_instruction = instruction[N - 1] && ~instruction[N - 2]; //es true si los bits más significativos son 10
    assign memoryInstruction = instruction[N - 1] && instruction[N -2]; //es true si los bits más significativos son 11

    // Outputs

    assign PcWriteEn = {
        instruction[N - 1] && ~instruction[N - 2] && ~instruction[N - 3] && instruction[N - 4], //1 si 1001
        instruction[N - 1] && ~instruction[N - 2] && ~instruction[N - 3] && ~instruction[N - 4], //1 si 1000
        instruction[N - 1] && instruction[N - 2] && instruction[N - 3] && instruction[N - 4] //1 si 1111
    };
	 


    assign MemoryWrite = memoryInstruction && ~instruction[N - 3] && ~instruction[N - 4];

    assign AluOpCode = instruction[N - 2:N - 4];

    assign preliminar_write_reg_from_1 = ~instruction[N - 1] & ~instruction[N - 2] & ~instruction[N - 3] & ~instruction[N - 4]; 
    assign WriteRegFrom[0] = preliminar_write_reg_from_1 ? 1'b0 : ~instruction[N - 1];
    assign WriteRegFrom[1] = (jump_instruction) ? jump_instruction : preliminar_write_reg_from_1;

    assign OverWriteNz = ~instruction[N - 1] & (|instruction[N - 2:N - 4]);

    assign RegToWrite = instruction[N - 5:N - 8];

	assign Immediate = instruction[N - 9:0]; 
    assign writeMemFrom = memoryInstruction && ~instruction[N - 3];

    assign regWriteEn = (memoryInstruction && instruction[N - 4]) | ~instruction[N -1];
    assign RegWriteEnSc = regWriteEn & (instruction[N - 6] || instruction[N - 5]);
    assign RegWriteEnVec = regWriteEn & ~instruction[N - 6] & ~instruction[N - 5];
	
endmodule