module top #(parameter N=8)(input clk, rst);
	
	processor proc(clk, rst);
	
endmodule