module key_expansion #(
    parameter regSize = 32,         // Size of each register (32 bits)
    parameter vecSize = 4           // Number of registers (4 words for AES-128)
)(
    input logic [vecSize-1:0][regSize-1:0] current_key, // Input key as a 2D array (4 x 32 bits)  
    input logic [vecSize-1:0][regSize-1:0] round,       // Round number as a 2D array
    output logic [vecSize-1:0][regSize-1:0] next_key    // Output next round key
);

    // Internal wire for the transformed word    
    logic [regSize-1:0] temp_word;    
    logic [regSize-1:0] sub_word_out; // Output from sub_word module  
    
    // Define round constants (Rcon) as a LUT    
    logic [31:0] rcon [0:10];     

    // Round constant initialization
    initial begin
        rcon[0] = 32'h01000000; rcon[1] = 32'h02000000;
        rcon[2] = 32'h04000000; rcon[3] = 32'h08000000;        
        rcon[4] = 32'h10000000; rcon[5] = 32'h20000000;
        rcon[6] = 32'h40000000; rcon[7] = 32'h80000000;        
        rcon[8] = 32'h1b000000; rcon[9] = 32'h36000000;
        rcon[10] = 32'h00000000; // Adjust as needed
    end
   
    // Define the S-box LUT
    logic [7:0] sbox [0:255]; // S-box for SubBytes transformation

    initial begin
		 sbox = '{
			  8'h63, 8'h7c, 8'h77, 8'h7b, 8'hf2, 8'h6b, 8'h6f, 8'hc5, 8'h30, 8'h01, 8'h67, 8'h2b, 8'hfe, 8'hd7, 8'hab, 8'h76,        
			  8'hca, 8'h82, 8'hc9, 8'h7d, 8'hfa, 8'h59, 8'h47, 8'hf0, 8'had, 8'hd4, 8'ha2, 8'haf, 8'h9c, 8'ha4, 8'h72, 8'hc0,
			  8'hb7, 8'hfd, 8'h93, 8'h26, 8'h36, 8'h3f, 8'hf7, 8'hcc, 8'h34, 8'ha5, 8'he5, 8'hf1, 8'h71, 8'hd8, 8'h31, 8'h15,        
			  8'h04, 8'hc7, 8'h23, 8'hc3, 8'h18, 8'h96, 8'h05, 8'h9a, 8'h07, 8'h12, 8'h80, 8'he2, 8'heb, 8'h27, 8'hb2, 8'h75,
			  8'h09, 8'h83, 8'h2c, 8'h1a, 8'h1b, 8'h6e, 8'h5a, 8'ha0, 8'h52, 8'h3b, 8'hd6, 8'hb3, 8'h29, 8'he3, 8'h2f, 8'h84,        
			  8'h53, 8'hd1, 8'h00, 8'hed, 8'h20, 8'hfc, 8'hb1, 8'h5b, 8'h6a, 8'hcb, 8'hbe, 8'h39, 8'h4a, 8'h4c, 8'h58, 8'hcf,
			  8'hd0, 8'hef, 8'haa, 8'hfb, 8'h43, 8'h4d, 8'h33, 8'h85, 8'h45, 8'hf9, 8'h02, 8'h7f, 8'h50, 8'h3c, 8'h9f, 8'ha8,        
			  8'h51, 8'ha3, 8'h40, 8'h8f, 8'h92, 8'h9d, 8'h38, 8'hf5, 8'hbc, 8'hb6, 8'hda, 8'h21, 8'h10, 8'hff, 8'hf3, 8'hd2,
			  8'hcd, 8'h0c, 8'h13, 8'hec, 8'h5f, 8'h97, 8'h44, 8'h17, 8'hc4, 8'ha7, 8'h7e, 8'h3d, 8'h64, 8'h5d, 8'h19, 8'h73,        
			  8'h60, 8'h81, 8'h4f, 8'hdc, 8'h22, 8'h2a, 8'h90, 8'h88, 8'h46, 8'hee, 8'hb8, 8'h14, 8'hde, 8'h5e, 8'h0b, 8'hdb,
			  8'he0, 8'h32, 8'h3a, 8'h0a, 8'h49, 8'h06, 8'h24, 8'h5c, 8'hc2, 8'hd3, 8'hac, 8'h62, 8'h91, 8'h95, 8'he4, 8'h79,        
			  8'he7, 8'hc8, 8'h37, 8'h6d, 8'h8d, 8'hd5, 8'h4e, 8'ha9, 8'h6c, 8'h56, 8'hf4, 8'hea, 8'h65, 8'h7a, 8'hae, 8'h08,
			  8'hba, 8'h78, 8'h25, 8'h2e, 8'h1c, 8'ha6, 8'hb4, 8'hc6, 8'he8, 8'hdd, 8'h74, 8'h1f, 8'h4b, 8'hbd, 8'h8b, 8'h8a,        
			  8'h70, 8'h3e, 8'hb5, 8'h66, 8'h48, 8'h03, 8'hf6, 8'h0e, 8'h61, 8'h35, 8'h57, 8'hb9, 8'h86, 8'hc1, 8'h1d, 8'h9e,
			  8'he1, 8'hf8, 8'h98, 8'h11, 8'h69, 8'hd9, 8'h8e, 8'h94, 8'h9b, 8'h1e, 8'h87, 8'he9, 8'hce, 8'h55, 8'h28, 8'hdf,        
			  8'h8c, 8'ha1, 8'h89, 8'h0d, 8'hbf, 8'he6, 8'h42, 8'h68, 8'h41, 8'h99, 8'h2d, 8'h0f, 8'hb0, 8'h54, 8'hbb, 8'h16
		 };
	  end

    // Substitution function using S-box
    function logic [regSize-1:0] sub_word(input logic [regSize-1:0] word_in);
        logic [regSize-1:0] word_out;
        begin
            word_out[31:24] = sbox[word_in[31:24]]; // SubBytes on each byte of the word
            word_out[23:16] = sbox[word_in[23:16]];
            word_out[15:8]  = sbox[word_in[15:8]];
            word_out[7:0]   = sbox[word_in[7:0]];
            return word_out;
        end
    endfunction
   
    // Compute the next key
    always_comb begin
        // Start with the last word of the current key        
        temp_word = current_key[vecSize-1];

        // Rotate the word left by 8 bits
        temp_word = {temp_word[23:0], temp_word[31:24]}; 

        // Apply the SubBytes (S-box) transformation
        temp_word = sub_word(temp_word);

        // XOR the result with the round constant for the current round
        // Use any element from the round 2D array (e.g., round[0][0])
        // Extract the least significant 4 bits of the round value (if needed)
        temp_word = temp_word ^ rcon[round[0][3:0]];

        // Generate the next key
        next_key[0] = current_key[0] ^ temp_word;        // XOR with the first word
        next_key[1] = current_key[1] ^ next_key[0];      // XOR with the previous result
        next_key[2] = current_key[2] ^ next_key[1];      // XOR with the previous result
        next_key[3] = current_key[3] ^ next_key[2];      // XOR with the previous result
    end
endmodule